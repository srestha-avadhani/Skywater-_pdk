magic
tech sky130A
timestamp 1640711282
<< nwell >>
rect 2885 1480 3070 1620
rect 3370 1480 4310 1620
rect -70 760 290 1460
rect 1395 1260 1995 1480
rect 1390 990 1995 1260
rect 2415 990 4310 1480
rect 1390 960 4310 990
rect 1800 460 1990 960
rect 2730 460 2780 960
rect 3370 955 4310 960
rect 3520 460 3570 955
<< locali >>
rect 1975 1355 1995 1585
rect 2565 1570 2585 1695
rect 3400 1645 3420 1780
rect 3370 1625 3420 1645
rect 2415 1550 2585 1570
rect 1435 1335 1995 1355
rect 1655 945 2060 965
rect 1655 905 1675 945
rect 2035 850 2060 945
rect 4330 410 4395 435
<< viali >>
rect 3400 1780 3420 1800
rect 3065 1675 3085 1695
rect 2870 1625 2890 1645
rect 2730 410 2750 430
rect 3520 410 3540 430
rect 1990 340 2010 360
rect 2780 340 2800 360
rect 3570 340 3590 360
<< metal1 >>
rect 3390 1805 3430 1810
rect 3390 1775 3395 1805
rect 3425 1775 3430 1805
rect 3390 1770 3430 1775
rect 2970 1710 3010 1715
rect 2970 1695 2975 1710
rect 2885 1680 2975 1695
rect 3005 1680 3010 1710
rect 2970 1675 3010 1680
rect 3055 1695 3095 1705
rect 3055 1675 3065 1695
rect 3085 1675 3095 1695
rect 3370 1680 4330 1695
rect 3055 1665 3095 1675
rect 2860 1650 2900 1655
rect 2860 1620 2865 1650
rect 2895 1620 2900 1650
rect 2860 1615 2900 1620
rect 3070 1525 3085 1665
rect 2415 1510 3085 1525
rect 2970 1355 3010 1360
rect 2970 1345 2975 1355
rect 2965 1330 2975 1345
rect 2970 1325 2975 1330
rect 3005 1335 3010 1355
rect 3005 1325 3490 1335
rect 2970 1320 3490 1325
rect 2730 595 2770 600
rect 2730 585 2735 595
rect 2685 570 2735 585
rect 1980 360 2020 370
rect 1980 340 1990 360
rect 2010 340 2020 360
rect 2685 340 2700 570
rect 2730 565 2735 570
rect 2765 565 2770 595
rect 2730 560 2770 565
rect 2720 435 2760 440
rect 2720 405 2725 435
rect 2755 405 2760 435
rect 2720 400 2760 405
rect 2765 360 2810 370
rect 2730 340 2750 355
rect 1980 330 2020 340
rect 1990 290 2005 330
rect 1955 275 2005 290
rect 1955 30 1970 275
rect 2735 30 2750 340
rect 2765 340 2780 360
rect 2800 340 2810 360
rect 3475 340 3490 1320
rect 3510 435 3550 440
rect 3510 405 3515 435
rect 3545 405 3550 435
rect 3510 400 3550 405
rect 3560 360 3600 370
rect 2765 330 2810 340
rect 2765 125 2780 330
rect 2765 110 2855 125
rect 1955 15 2750 30
rect 2840 30 2855 110
rect 3530 30 3545 355
rect 3560 340 3570 360
rect 3590 340 3600 360
rect 3560 330 3600 340
rect 3575 140 3590 330
rect 3575 125 3650 140
rect 2840 15 3545 30
rect 3635 30 3650 125
rect 4315 30 4330 1680
rect 3635 15 4330 30
<< via1 >>
rect 3395 1800 3425 1805
rect 3395 1780 3400 1800
rect 3400 1780 3420 1800
rect 3420 1780 3425 1800
rect 3395 1775 3425 1780
rect 2975 1680 3005 1710
rect 2865 1645 2895 1650
rect 2865 1625 2870 1645
rect 2870 1625 2890 1645
rect 2890 1625 2895 1645
rect 2865 1620 2895 1625
rect 2975 1325 3005 1355
rect 2735 565 2765 595
rect 2725 430 2755 435
rect 2725 410 2730 430
rect 2730 410 2750 430
rect 2750 410 2755 430
rect 2725 405 2755 410
rect 3515 430 3545 435
rect 3515 410 3520 430
rect 3520 410 3540 430
rect 3540 410 3545 430
rect 3515 405 3545 410
<< metal2 >>
rect 3385 1805 3435 1820
rect -185 1790 3395 1805
rect 3385 1775 3395 1790
rect 3425 1775 3435 1805
rect 3385 1765 3435 1775
rect 2965 1710 3015 1720
rect 2965 1680 2975 1710
rect 3005 1680 3015 1710
rect 2965 1670 3015 1680
rect 2855 1650 2905 1660
rect 2855 1620 2865 1650
rect 2895 1645 2905 1650
rect 2895 1620 2915 1645
rect 2855 1610 2915 1620
rect 2900 995 2915 1610
rect 2985 1365 3000 1670
rect 2965 1355 3015 1365
rect 2965 1325 2975 1355
rect 3005 1325 3015 1355
rect 2965 1315 3015 1325
rect 2745 980 2915 995
rect 2745 605 2760 980
rect 2725 595 2775 605
rect 2725 565 2735 595
rect 2765 565 2775 595
rect 2725 555 2775 565
rect -185 430 -155 450
rect 1955 430 1990 450
rect 2735 445 2780 450
rect 3520 445 3570 450
rect 2715 435 2780 445
rect 1955 340 1970 430
rect 2715 405 2725 435
rect 2755 430 2780 435
rect 3505 435 3570 445
rect 2755 405 2765 430
rect 2715 395 2765 405
rect 3505 405 3515 435
rect 3545 430 3570 435
rect 3545 405 3555 430
rect 3505 395 3555 405
<< metal4 >>
rect 1885 1850 2040 1885
rect 2345 1865 2590 1895
rect 2885 1865 3070 1895
rect 1885 1530 1915 1850
rect 2350 1080 2785 1110
rect 2885 1080 3070 1110
rect 1995 960 2415 995
rect 2725 930 2815 960
rect 3515 930 3605 960
rect 1915 15 2005 45
rect 2715 15 2810 45
rect 3510 15 3600 45
use tspc  tspc_2
timestamp 1640710665
transform 1 0 3640 0 1 495
box -70 -565 690 465
use tspc  tspc_1
timestamp 1640710665
transform 1 0 2850 0 1 495
box -70 -565 690 465
use tspc  tspc_0
timestamp 1640710665
transform 1 0 2060 0 1 495
box -70 -565 690 465
use prescaler  prescaler_0
timestamp 1640711282
transform 1 0 25 0 1 200
box -210 -270 1930 1790
use and  and_0
timestamp 1640698682
transform -1 0 2330 0 -1 1465
box -85 -490 335 475
use nor  nor_0
timestamp 1640700690
transform -1 0 2830 0 -1 1605
box -55 -300 290 610
use nor  nor_1
timestamp 1640700690
transform -1 0 3315 0 -1 1605
box -55 -300 290 610
<< labels >>
rlabel metal4 1915 15 2005 45 1 gnd
rlabel metal4 2715 15 2810 45 1 gnd
rlabel space 3510 15 3605 45 1 gnd
rlabel space 3515 930 3610 960 1 vdd
rlabel metal4 2725 930 2815 960 1 vdd
rlabel metal4 1995 965 2415 995 1 vdd
rlabel metal4 2350 1080 2585 1110 1 vdd
rlabel metal4 2885 1080 3070 1110 1 vdd
rlabel metal4 1885 1560 1915 1885 1 gnd
rlabel metal4 1915 1850 2035 1885 1 gnd
rlabel locali 4330 410 4395 435 1 Out
rlabel metal2 -185 430 -155 450 1 clk
rlabel metal2 -185 1790 225 1805 1 mc2
<< end >>
