* SPICE3 file created from divider.ext - technology: sky130A
.lib "/home/sresthavadhani/sky/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param SUPPLY = 1.8
.global vdd gnd

Vdd vdd gnd 'SUPPLY'
Vin_clk clk gnd pulse 0 1.8 0 0 0 1n 2n
Vin_mc mc2 gnd 1.8


X0 and_0/A nor_0/B gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 and_0/A nor_0/A gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 nor_0/Z1 nor_0/A vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=150000u
X3 and_0/A nor_0/B nor_0/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=150000u
X4 and_0/B nor_1/B gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 and_0/B mc2 gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 nor_1/Z1 mc2 vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=150000u
X7 and_0/B nor_1/B nor_1/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=150000u
X8 prescaler_0/tspc_0/Z3 prescaler_0/tspc_0/Z2 prescaler_0/tspc_0/Z4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X9 prescaler_0/tspc_0/Z4 clk gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X10 prescaler_0/tspc_0/Z1 prescaler_0/tspc_0/D vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X11 prescaler_0/tspc_0/Z2 prescaler_0/tspc_0/D gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X12 prescaler_0/Out prescaler_0/tspc_0/a_740_n680# vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X13 prescaler_0/tspc_0/a_740_n680# prescaler_0/tspc_0/Z3 vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X14 prescaler_0/tspc_0/Z2 clk prescaler_0/tspc_0/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X15 prescaler_0/Out prescaler_0/tspc_0/a_740_n680# gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X16 prescaler_0/tspc_0/a_740_n680# clk prescaler_0/tspc_0/a_630_n680# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 prescaler_0/tspc_0/a_630_n680# prescaler_0/tspc_0/Z3 gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 prescaler_0/tspc_0/Z3 clk vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X19 prescaler_0/tspc_1/Z3 prescaler_0/tspc_1/Z2 prescaler_0/tspc_1/Z4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X20 prescaler_0/tspc_1/Z4 clk gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X21 prescaler_0/tspc_1/Z1 prescaler_0/Out vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X22 prescaler_0/tspc_1/Z2 prescaler_0/Out gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X23 prescaler_0/tspc_1/Q prescaler_0/m1_2700_2190# vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X24 prescaler_0/m1_2700_2190# prescaler_0/tspc_1/Z3 vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X25 prescaler_0/tspc_1/Z2 clk prescaler_0/tspc_1/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X26 prescaler_0/tspc_1/Q prescaler_0/m1_2700_2190# gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X27 prescaler_0/m1_2700_2190# clk prescaler_0/tspc_1/a_630_n680# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 prescaler_0/tspc_1/a_630_n680# prescaler_0/tspc_1/Z3 gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 prescaler_0/tspc_1/Z3 clk vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X30 prescaler_0/tspc_2/Z3 prescaler_0/tspc_2/Z2 prescaler_0/tspc_2/Z4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X31 prescaler_0/tspc_2/Z4 clk gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X32 prescaler_0/tspc_2/Z1 prescaler_0/tspc_2/D vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X33 prescaler_0/tspc_2/Z2 prescaler_0/tspc_2/D gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X34 prescaler_0/tspc_2/Q prescaler_0/tspc_2/a_740_n680# vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X35 prescaler_0/tspc_2/a_740_n680# prescaler_0/tspc_2/Z3 vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X36 prescaler_0/tspc_2/Z2 clk prescaler_0/tspc_2/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X37 prescaler_0/tspc_2/Q prescaler_0/tspc_2/a_740_n680# gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X38 prescaler_0/tspc_2/a_740_n680# clk prescaler_0/tspc_2/a_630_n680# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 prescaler_0/tspc_2/a_630_n680# prescaler_0/tspc_2/Z3 gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 prescaler_0/tspc_2/Z3 clk vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X41 prescaler_0/tspc_0/D prescaler_0/tspc_2/Q vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X42 prescaler_0/tspc_0/D prescaler_0/tspc_1/Q vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X43 prescaler_0/nand_0/z1 prescaler_0/tspc_2/Q gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 prescaler_0/tspc_0/D prescaler_0/tspc_1/Q prescaler_0/nand_0/z1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 prescaler_0/tspc_2/D and_0/OUT vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X46 prescaler_0/tspc_2/D prescaler_0/m1_2700_2190# vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X47 prescaler_0/nand_1/z1 and_0/OUT gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 prescaler_0/tspc_2/D prescaler_0/m1_2700_2190# prescaler_0/nand_1/z1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X49 tspc_0/Z3 tspc_0/Z2 tspc_0/Z4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X50 tspc_0/Z4 prescaler_0/Out gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X51 tspc_0/Z1 nor_0/A vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X52 tspc_0/Z2 nor_0/A gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X53 tspc_0/Q nor_0/A vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X54 nor_0/A tspc_0/Z3 vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X55 tspc_0/Z2 prescaler_0/Out tspc_0/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X56 tspc_0/Q nor_0/A gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X57 nor_0/A prescaler_0/Out tspc_0/a_630_n680# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 tspc_0/a_630_n680# tspc_0/Z3 gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 tspc_0/Z3 prescaler_0/Out vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X60 tspc_1/Z3 tspc_1/Z2 tspc_1/Z4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X61 tspc_1/Z4 tspc_0/Q gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X62 tspc_1/Z1 nor_0/B vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X63 tspc_1/Z2 nor_0/B gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X64 tspc_1/Q nor_0/B vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X65 nor_0/B tspc_1/Z3 vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X66 tspc_1/Z2 tspc_0/Q tspc_1/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X67 tspc_1/Q nor_0/B gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X68 nor_0/B tspc_0/Q tspc_1/a_630_n680# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X69 tspc_1/a_630_n680# tspc_1/Z3 gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X70 tspc_1/Z3 tspc_0/Q vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X71 tspc_2/Z3 tspc_2/Z2 tspc_2/Z4 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X72 tspc_2/Z4 tspc_1/Q gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.8e+06u l=150000u
X73 tspc_2/Z1 nor_1/B vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X74 tspc_2/Z2 nor_1/B gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=450000u l=150000u
X75 Out nor_1/B vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=4e+06u l=150000u
X76 nor_1/B tspc_2/Z3 vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X77 tspc_2/Z2 tspc_1/Q tspc_2/Z1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.8e+06u l=150000u
X78 Out nor_1/B gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X79 nor_1/B tspc_1/Q tspc_2/a_630_n680# VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X80 tspc_2/a_630_n680# tspc_2/Z3 gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X81 tspc_2/Z3 tspc_1/Q vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.9e+06u l=150000u
X82 and_0/OUT and_0/out1 vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=3.8e+06u l=150000u
X83 and_0/Z1 and_0/A gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X84 and_0/out1 and_0/A vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.6e+06u l=150000u
X85 and_0/out1 and_0/B and_0/Z1 VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2e+06u l=150000u
X86 and_0/OUT and_0/out1 gnd VSUBS sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=150000u
X87 and_0/out1 and_0/B vdd VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.6e+06u l=150000u
C0 prescaler_0/tspc_2/Z2 clk 0.11fF
C1 gnd prescaler_0/tspc_1/Q 0.83fF
C2 mc2 and_0/OUT 0.05fF
C3 prescaler_0/tspc_1/Z4 vdd 0.01fF
C4 gnd prescaler_0/tspc_2/Z4 0.44fF
C5 clk prescaler_0/tspc_2/Q 0.05fF
C6 nor_0/A tspc_0/Z2 0.23fF
C7 nor_0/B tspc_1/Z3 0.38fF
C8 prescaler_0/tspc_0/Z2 prescaler_0/tspc_0/Z1 1.07fF
C9 gnd prescaler_0/tspc_2/Z2 0.16fF
C10 vdd and_0/out1 1.44fF
C11 prescaler_0/tspc_1/Q prescaler_0/nand_0/z1 0.22fF
C12 gnd prescaler_0/tspc_2/Q 0.35fF
C13 and_0/OUT and_0/Z1 0.04fF
C14 vdd clk 0.27fF
C15 nor_0/A tspc_1/Z2 0.15fF
C16 nor_0/A prescaler_0/tspc_1/Q 0.03fF
C17 gnd prescaler_0/tspc_1/a_630_n680# 0.00fF
C18 prescaler_0/nand_1/z1 and_0/OUT 0.01fF
C19 gnd tspc_2/Z4 0.44fF
C20 prescaler_0/tspc_1/Z1 vdd 0.58fF
C21 vdd tspc_1/Z1 0.01fF
C22 vdd gnd 0.26fF
C23 nor_1/B Out 0.22fF
C24 gnd prescaler_0/tspc_2/D 0.14fF
C25 tspc_2/Z2 tspc_2/Z4 0.36fF
C26 tspc_2/Z4 tspc_2/a_630_n680# 0.12fF
C27 prescaler_0/tspc_2/Q prescaler_0/nand_0/z1 0.01fF
C28 prescaler_0/Out prescaler_0/tspc_1/Z2 0.19fF
C29 gnd nor_1/Z1 0.01fF
C30 vdd tspc_2/Z2 0.36fF
C31 gnd tspc_0/Z4 0.00fF
C32 clk prescaler_0/tspc_2/Z3 0.45fF
C33 prescaler_0/tspc_2/a_630_n680# clk 0.01fF
C34 prescaler_0/tspc_0/Z3 prescaler_0/tspc_0/D 0.05fF
C35 prescaler_0/Out tspc_0/Z3 0.45fF
C36 vdd prescaler_0/nand_0/z1 0.01fF
C37 tspc_0/Q tspc_0/Z3 0.05fF
C38 tspc_2/Z1 tspc_2/Z2 1.07fF
C39 and_0/B and_0/A 0.18fF
C40 gnd prescaler_0/tspc_2/Z3 0.27fF
C41 vdd nor_0/A 0.83fF
C42 prescaler_0/tspc_2/Z2 and_0/OUT 0.05fF
C43 prescaler_0/tspc_2/a_630_n680# gnd 0.61fF
C44 tspc_0/Q tspc_1/Z4 0.15fF
C45 prescaler_0/tspc_1/Z4 prescaler_0/Out 0.28fF
C46 prescaler_0/tspc_2/Q and_0/OUT 0.04fF
C47 prescaler_0/tspc_0/a_630_n680# prescaler_0/Out 0.04fF
C48 prescaler_0/tspc_0/D prescaler_0/tspc_1/Q 0.32fF
C49 and_0/A nor_0/B 0.26fF
C50 clk prescaler_0/Out 0.51fF
C51 prescaler_0/tspc_1/a_630_n680# prescaler_0/m1_2700_2190# 0.19fF
C52 vdd and_0/OUT 1.59fF
C53 gnd tspc_1/Q 0.33fF
C54 prescaler_0/tspc_2/Q prescaler_0/tspc_0/D 0.04fF
C55 and_0/A gnd 0.09fF
C56 tspc_1/Q tspc_2/a_630_n680# 0.01fF
C57 tspc_1/Q tspc_2/Z2 0.14fF
C58 prescaler_0/tspc_2/D prescaler_0/m1_2700_2190# 0.16fF
C59 tspc_1/Z1 tspc_1/Z4 0.00fF
C60 prescaler_0/tspc_1/Z1 prescaler_0/Out 0.08fF
C61 gnd prescaler_0/Out 0.46fF
C62 gnd nor_1/B 0.96fF
C63 tspc_0/a_630_n680# tspc_0/Z2 0.01fF
C64 gnd tspc_0/Q 0.33fF
C65 nor_1/B tspc_2/Z2 0.40fF
C66 nor_1/B tspc_2/a_630_n680# 0.35fF
C67 vdd prescaler_0/tspc_0/D 0.90fF
C68 prescaler_0/tspc_0/Z2 prescaler_0/tspc_0/Z4 0.36fF
C69 prescaler_0/tspc_1/Z3 prescaler_0/tspc_1/Q 0.21fF
C70 and_0/B and_0/out1 0.18fF
C71 nor_0/B tspc_1/Z4 0.21fF
C72 vdd prescaler_0/tspc_2/D 0.07fF
C73 clk prescaler_0/tspc_2/a_740_n680# 0.01fF
C74 mc2 and_0/Z1 0.09fF
C75 prescaler_0/tspc_0/a_630_n680# prescaler_0/tspc_0/Z4 0.12fF
C76 prescaler_0/tspc_0/a_740_n680# prescaler_0/tspc_0/Z3 0.33fF
C77 nor_0/A prescaler_0/Out 0.15fF
C78 prescaler_0/tspc_0/D prescaler_0/tspc_0/Z1 0.03fF
C79 gnd tspc_1/Z4 0.00fF
C80 and_0/B gnd 0.45fF
C81 nor_0/A tspc_0/Q 0.55fF
C82 prescaler_0/tspc_1/Z4 gnd 0.00fF
C83 gnd prescaler_0/tspc_2/a_740_n680# 0.22fF
C84 prescaler_0/tspc_0/a_630_n680# gnd 0.00fF
C85 prescaler_0/tspc_2/Z1 prescaler_0/tspc_2/Z4 0.00fF
C86 clk prescaler_0/tspc_0/Z4 0.12fF
C87 tspc_2/Z3 Out 0.05fF
C88 prescaler_0/tspc_0/a_740_n680# prescaler_0/tspc_1/Q 0.15fF
C89 prescaler_0/tspc_2/Z1 prescaler_0/tspc_2/Z2 1.07fF
C90 prescaler_0/tspc_1/a_630_n680# prescaler_0/tspc_1/Z2 0.01fF
C91 tspc_0/Z4 tspc_0/Z1 0.00fF
C92 vdd prescaler_0/tspc_1/Z3 0.67fF
C93 gnd prescaler_0/tspc_0/Z4 0.44fF
C94 gnd nor_0/B 0.99fF
C95 and_0/B nor_0/A 0.08fF
C96 nor_0/B tspc_2/Z2 0.20fF
C97 gnd gnd 0.07fF
C98 tspc_1/Z3 tspc_1/Z4 0.65fF
C99 prescaler_0/tspc_2/Z2 mc2 0.24fF
C100 vdd prescaler_0/tspc_2/Z1 0.58fF
C101 gnd tspc_2/a_630_n680# 0.00fF
C102 vdd tspc_0/Z1 0.01fF
C103 tspc_0/Z4 tspc_0/Z3 0.65fF
C104 prescaler_0/tspc_1/Z4 prescaler_0/tspc_1/a_630_n680# 0.12fF
C105 vdd prescaler_0/tspc_0/a_740_n680# 0.52fF
C106 nor_0/A nor_0/B 1.22fF
C107 and_0/B and_0/OUT 0.01fF
C108 gnd prescaler_0/nand_0/z1 0.01fF
C109 prescaler_0/tspc_0/Z3 prescaler_0/tspc_1/Q 0.13fF
C110 prescaler_0/tspc_1/Z4 prescaler_0/m1_2700_2190# 0.08fF
C111 vdd mc2 0.06fF
C112 tspc_1/a_630_n680# tspc_1/Z2 0.01fF
C113 clk prescaler_0/tspc_1/a_630_n680# 0.01fF
C114 prescaler_0/tspc_2/Z1 prescaler_0/tspc_2/Z3 0.06fF
C115 clk prescaler_0/tspc_2/D 0.26fF
C116 gnd tspc_1/Z3 0.27fF
C117 clk prescaler_0/m1_2700_2190# 0.01fF
C118 gnd prescaler_0/tspc_1/a_630_n680# 0.61fF
C119 vdd and_0/Z1 0.01fF
C120 gnd tspc_2/Z3 0.27fF
C121 tspc_2/Z3 tspc_2/Z2 0.16fF
C122 prescaler_0/tspc_1/Z3 prescaler_0/Out 0.11fF
C123 tspc_2/Z3 tspc_2/a_630_n680# 0.05fF
C124 gnd prescaler_0/tspc_2/D 0.05fF
C125 vdd prescaler_0/nand_1/z1 0.01fF
C126 vdd prescaler_0/tspc_0/Z3 0.67fF
C127 vdd tspc_0/Z2 0.37fF
C128 prescaler_0/Out tspc_0/a_630_n680# 0.01fF
C129 prescaler_0/tspc_2/a_630_n680# mc2 0.19fF
C130 prescaler_0/tspc_2/Z2 prescaler_0/tspc_2/Z4 0.36fF
C131 gnd prescaler_0/m1_2700_2190# 0.22fF
C132 gnd tspc_0/Z4 0.44fF
C133 prescaler_0/tspc_2/Q prescaler_0/tspc_1/Q 0.19fF
C134 tspc_0/Z3 tspc_0/Z1 0.06fF
C135 tspc_0/Q tspc_0/a_630_n680# 0.04fF
C136 prescaler_0/tspc_0/Z4 prescaler_0/tspc_0/D 0.11fF
C137 vdd and_0/out1 0.01fF
C138 vdd nor_0/Z1 0.75fF
C139 vdd tspc_1/Z2 0.36fF
C140 prescaler_0/tspc_0/Z3 prescaler_0/tspc_0/Z1 0.06fF
C141 gnd prescaler_0/tspc_0/D 0.04fF
C142 vdd prescaler_0/tspc_1/Q 0.64fF
C143 vdd prescaler_0/tspc_2/Z4 0.01fF
C144 prescaler_0/tspc_1/Z1 vdd 0.01fF
C145 prescaler_0/Out prescaler_0/tspc_0/a_740_n680# 0.21fF
C146 nor_0/A prescaler_0/m1_2700_2190# 0.01fF
C147 nor_0/A tspc_0/Z4 0.21fF
C148 vdd prescaler_0/tspc_2/Z2 0.37fF
C149 prescaler_0/tspc_1/Z4 prescaler_0/tspc_1/Z2 0.36fF
C150 and_0/A and_0/out1 0.01fF
C151 mc2 nor_1/B 0.15fF
C152 vdd prescaler_0/tspc_2/Q 0.70fF
C153 and_0/OUT prescaler_0/tspc_2/D 0.03fF
C154 prescaler_0/tspc_2/Z3 prescaler_0/tspc_2/Z4 0.65fF
C155 vdd tspc_2/Z4 0.01fF
C156 clk prescaler_0/tspc_1/Z2 0.11fF
C157 and_0/A gnd 0.53fF
C158 and_0/OUT prescaler_0/m1_2700_2190# 0.14fF
C159 nor_0/B tspc_0/a_630_n680# 0.01fF
C160 prescaler_0/tspc_2/a_630_n680# prescaler_0/tspc_2/Z4 0.12fF
C161 prescaler_0/tspc_0/Z2 prescaler_0/tspc_0/a_630_n680# 0.01fF
C162 prescaler_0/tspc_2/Z2 prescaler_0/tspc_2/Z3 0.16fF
C163 vdd nor_1/Z1 0.75fF
C164 gnd Out 0.29fF
C165 prescaler_0/Out tspc_0/Z2 0.11fF
C166 prescaler_0/Out prescaler_0/tspc_0/Z3 0.05fF
C167 prescaler_0/tspc_2/a_630_n680# prescaler_0/tspc_2/Z2 0.01fF
C168 prescaler_0/tspc_2/Q prescaler_0/tspc_2/Z3 0.05fF
C169 prescaler_0/tspc_1/Z1 prescaler_0/tspc_1/Z2 1.07fF
C170 gnd prescaler_0/tspc_1/Z2 0.17fF
C171 gnd tspc_0/a_630_n680# 0.00fF
C172 tspc_1/Q tspc_1/a_630_n680# 0.04fF
C173 and_0/B mc2 0.20fF
C174 tspc_2/a_630_n680# Out 0.04fF
C175 tspc_2/Z1 tspc_2/Z4 0.00fF
C176 prescaler_0/tspc_2/a_630_n680# prescaler_0/tspc_2/Q 0.04fF
C177 prescaler_0/tspc_0/Z2 clk 0.11fF
C178 vdd tspc_2/Z1 0.58fF
C179 vdd prescaler_0/tspc_0/Z1 0.58fF
C180 vdd and_0/OUT 0.01fF
C181 gnd tspc_0/Z3 0.27fF
C182 nor_0/A tspc_0/Z1 0.03fF
C183 tspc_1/a_630_n680# nor_1/B 0.00fF
C184 prescaler_0/tspc_1/Z4 clk 0.12fF
C185 prescaler_0/tspc_0/a_740_n680# prescaler_0/tspc_0/Z4 0.08fF
C186 and_0/A nor_0/A 0.01fF
C187 vdd prescaler_0/tspc_2/Z3 0.67fF
C188 prescaler_0/tspc_0/a_630_n680# clk 0.01fF
C189 tspc_0/Q tspc_1/Z2 0.14fF
C190 tspc_1/a_630_n680# tspc_0/Q 0.01fF
C191 prescaler_0/Out prescaler_0/tspc_1/Q 0.91fF
C192 prescaler_0/tspc_0/Z2 gnd 0.16fF
C193 and_0/B and_0/Z1 0.07fF
C194 gnd tspc_1/Z4 0.44fF
C195 mc2 nor_0/B 0.07fF
C196 prescaler_0/tspc_1/Z4 prescaler_0/tspc_1/Z1 0.00fF
C197 prescaler_0/tspc_1/Z4 gnd 0.44fF
C198 prescaler_0/tspc_0/a_630_n680# gnd 0.63fF
C199 vdd prescaler_0/tspc_0/D 0.06fF
C200 gnd mc2 0.13fF
C201 prescaler_0/tspc_1/Z3 prescaler_0/tspc_1/a_630_n680# 0.05fF
C202 tspc_1/Q tspc_2/Z4 0.15fF
C203 nor_0/A tspc_0/Z3 0.38fF
C204 and_0/B nor_0/Z1 0.18fF
C205 gnd and_0/out1 0.23fF
C206 vdd tspc_1/Q 0.72fF
C207 gnd clk 0.07fF
C208 prescaler_0/tspc_2/a_630_n680# prescaler_0/tspc_2/Z3 0.05fF
C209 tspc_1/Z1 tspc_1/Z2 1.07fF
C210 nor_0/A tspc_1/Z4 0.02fF
C211 nor_1/B tspc_2/Z4 0.22fF
C212 and_0/OUT prescaler_0/tspc_1/Z2 0.06fF
C213 prescaler_0/tspc_1/Z3 prescaler_0/m1_2700_2190# 0.33fF
C214 prescaler_0/tspc_0/Z3 prescaler_0/tspc_0/Z4 0.65fF
C215 gnd and_0/Z1 0.02fF
C216 vdd prescaler_0/Out 0.75fF
C217 vdd nor_1/B 0.55fF
C218 tspc_0/Z4 tspc_0/a_630_n680# 0.12fF
C219 prescaler_0/tspc_2/a_740_n680# prescaler_0/tspc_2/Z4 0.08fF
C220 vdd tspc_0/Q 0.72fF
C221 nor_1/B nor_1/Z1 0.06fF
C222 tspc_2/Z1 tspc_1/Q 0.01fF
C223 gnd prescaler_0/nand_1/z1 0.01fF
C224 nor_0/B nor_0/Z1 0.06fF
C225 gnd tspc_2/Z2 0.16fF
C226 prescaler_0/tspc_2/Z1 prescaler_0/tspc_2/D 0.15fF
C227 gnd tspc_2/a_630_n680# 0.61fF
C228 nor_0/B tspc_1/Z2 0.30fF
C229 tspc_1/a_630_n680# nor_0/B 0.35fF
C230 prescaler_0/tspc_0/Z2 and_0/OUT 0.06fF
C231 tspc_2/Z2 tspc_2/a_630_n680# 0.01fF
C232 prescaler_0/tspc_0/Z4 prescaler_0/tspc_1/Q 0.21fF
C233 tspc_2/Z1 nor_1/B 0.03fF
C234 prescaler_0/tspc_2/Q prescaler_0/tspc_2/a_740_n680# 0.20fF
C235 gnd prescaler_0/nand_0/z1 0.16fF
C236 gnd tspc_1/a_630_n680# 0.00fF
C237 and_0/B vdd 0.20fF
C238 nor_0/A gnd 0.90fF
C239 gnd prescaler_0/tspc_2/Z4 0.00fF
C240 vdd tspc_1/Z1 0.58fF
C241 vdd prescaler_0/tspc_2/a_740_n680# 0.52fF
C242 and_0/B nor_1/Z1 0.78fF
C243 prescaler_0/tspc_0/Z2 prescaler_0/tspc_0/D 0.09fF
C244 and_0/OUT and_0/out1 0.31fF
C245 vdd prescaler_0/tspc_2/Z1 0.02fF
C246 clk and_0/OUT 0.04fF
C247 nor_0/B tspc_2/Z4 0.02fF
C248 tspc_1/Q nor_1/B 0.22fF
C249 vdd prescaler_0/tspc_0/Z4 0.01fF
C250 vdd nor_0/B 0.30fF
C251 gnd and_0/OUT 0.26fF
C252 nor_0/B nor_1/Z1 0.26fF
C253 prescaler_0/nand_1/z1 prescaler_0/tspc_2/D 0.24fF
C254 prescaler_0/tspc_1/Z3 prescaler_0/tspc_1/Z2 0.16fF
C255 gnd tspc_2/Z4 0.00fF
C256 prescaler_0/tspc_2/a_740_n680# prescaler_0/tspc_2/Z3 0.33fF
C257 tspc_1/Z3 tspc_1/Z2 0.16fF
C258 tspc_1/a_630_n680# tspc_1/Z3 0.05fF
C259 clk prescaler_0/tspc_0/D 0.29fF
C260 prescaler_0/nand_1/z1 prescaler_0/m1_2700_2190# 0.07fF
C261 prescaler_0/tspc_2/a_630_n680# prescaler_0/tspc_2/a_740_n680# 0.19fF
C262 tspc_0/Z4 tspc_0/Z2 0.36fF
C263 prescaler_0/tspc_0/Z4 prescaler_0/tspc_0/Z1 0.00fF
C264 prescaler_0/tspc_1/a_630_n680# prescaler_0/tspc_1/Q 0.04fF
C265 gnd prescaler_0/tspc_0/D 0.05fF
C266 tspc_0/a_630_n680# tspc_0/Z3 0.05fF
C267 prescaler_0/tspc_2/Z4 prescaler_0/tspc_2/D 0.11fF
C268 prescaler_0/tspc_1/Q prescaler_0/m1_2700_2190# 0.38fF
C269 and_0/A mc2 0.16fF
C270 prescaler_0/tspc_1/Z4 prescaler_0/tspc_1/Z3 0.65fF
C271 prescaler_0/tspc_0/a_740_n680# prescaler_0/tspc_1/Z2 0.01fF
C272 prescaler_0/tspc_2/Z2 prescaler_0/tspc_2/D 0.09fF
C273 prescaler_0/tspc_2/a_630_n680# gnd 0.00fF
C274 prescaler_0/tspc_0/D prescaler_0/nand_0/z1 0.21fF
C275 and_0/B nor_1/B 0.29fF
C276 vdd nor_0/Z1 0.02fF
C277 vdd tspc_1/Z3 0.67fF
C278 tspc_0/Q tspc_1/Z1 0.01fF
C279 tspc_2/Z3 tspc_2/Z4 0.65fF
C280 prescaler_0/tspc_1/Z3 clk 0.45fF
C281 tspc_1/Q nor_0/B 0.51fF
C282 vdd tspc_2/Z3 0.67fF
C283 tspc_0/Z2 tspc_0/Z1 1.07fF
C284 vdd prescaler_0/tspc_2/D 1.18fF
C285 nor_0/B nor_1/B 0.48fF
C286 prescaler_0/tspc_1/Z4 prescaler_0/tspc_0/a_740_n680# 0.01fF
C287 prescaler_0/tspc_1/Z1 prescaler_0/tspc_1/Z3 0.06fF
C288 prescaler_0/tspc_1/Z3 gnd 0.27fF
C289 vdd prescaler_0/m1_2700_2190# 0.59fF
C290 prescaler_0/tspc_0/a_630_n680# prescaler_0/tspc_0/a_740_n680# 0.19fF
C291 vdd tspc_0/Z4 0.01fF
C292 tspc_0/Q nor_0/B 0.22fF
C293 tspc_2/Z1 tspc_2/Z3 0.06fF
C294 gnd tspc_0/a_630_n680# 0.62fF
C295 and_0/A nor_0/Z1 0.80fF
C296 clk prescaler_0/tspc_0/a_740_n680# 0.14fF
C297 prescaler_0/tspc_2/Z3 prescaler_0/tspc_2/D 0.05fF
C298 tspc_0/Z2 tspc_0/Z3 0.16fF
C299 mc2 and_0/out1 0.06fF
C300 vdd vdd 0.23fF
C301 prescaler_0/tspc_0/Z2 prescaler_0/tspc_0/Z3 0.16fF
C302 prescaler_0/tspc_1/Z2 prescaler_0/tspc_1/Q 0.06fF
C303 vdd nor_1/Z1 0.02fF
C304 and_0/B nor_0/B 0.35fF
C305 gnd prescaler_0/tspc_0/a_740_n680# 0.22fF
C306 nor_0/B tspc_1/Z1 0.03fF
C307 nor_0/A tspc_0/a_630_n680# 0.35fF
C308 tspc_1/Q tspc_1/Z3 0.05fF
C309 prescaler_0/tspc_0/a_630_n680# prescaler_0/tspc_0/Z3 0.05fF
C310 gnd mc2 1.02fF
C311 tspc_1/Q tspc_2/Z3 0.45fF
C312 and_0/out1 and_0/Z1 0.36fF
C313 and_0/B gnd 0.08fF
C314 vdd prescaler_0/tspc_0/Z1 0.02fF
C315 vdd tspc_2/Z1 0.01fF
C316 tspc_1/Z2 tspc_1/Z4 0.36fF
C317 tspc_1/a_630_n680# tspc_1/Z4 0.12fF
C318 prescaler_0/tspc_0/Z2 prescaler_0/tspc_1/Q 0.06fF
C319 vdd tspc_0/Z1 0.58fF
C320 and_0/A vdd 0.11fF
C321 tspc_2/Z3 nor_1/B 0.38fF
C322 tspc_0/Q tspc_1/Z3 0.45fF
C323 clk prescaler_0/tspc_0/Z3 0.64fF
C324 prescaler_0/tspc_1/Z4 prescaler_0/tspc_1/Q 0.16fF
C325 gnd and_0/Z1 0.41fF
C326 vdd Out 0.61fF
C327 gnd prescaler_0/tspc_0/Z4 0.02fF
C328 vdd prescaler_0/tspc_1/Z2 0.38fF
C329 prescaler_0/Out prescaler_0/m1_2700_2190# 0.11fF
C330 gnd prescaler_0/nand_1/z1 0.16fF
C331 prescaler_0/Out tspc_0/Z4 0.12fF
C332 nor_0/A mc2 0.04fF
C333 gnd prescaler_0/tspc_0/Z3 0.27fF
C334 gnd tspc_0/Z2 0.16fF
C335 clk prescaler_0/tspc_1/Q 0.60fF
C336 vdd tspc_0/Z3 0.67fF
C337 clk prescaler_0/tspc_2/Z4 0.12fF
C338 gnd nor_0/Z1 0.01fF
C339 tspc_1/Z3 tspc_1/Z1 0.06fF
C340 gnd tspc_1/Z2 0.16fF
C341 gnd tspc_1/a_630_n680# 0.62fF
C342 prescaler_0/tspc_0/Z2 vdd 0.37fF
C343 vdd tspc_1/Z4 0.01fF
C344 and_0/Z1 VDD 0.31fF 
C345 and_0/B VDD 1.98fF 
C346 and_0/A VDD 1.56fF 
C347 and_0/out1 VDD 1.26fF 
C348 gnd VDD 1.57fF
C349 vdd VDD 1.47fF
C350 tspc_2/a_630_n680# VDD 0.52fF 
C351 tspc_2/Z4 VDD 0.41fF 
C352 Out VDD 0.70fF 
C353 tspc_2/Z3 VDD 1.33fF 
C354 tspc_2/Z2 VDD 0.91fF 
C355 tspc_2/Z1 VDD 0.41fF 
C356 tspc_1/Q VDD 1.46fF 
C357 nor_1/B VDD 5.20fF 
C358 tspc_1/a_630_n680# VDD 0.52fF 
C359 tspc_1/Z4 VDD 0.41fF 
C360 tspc_1/Z3 VDD 1.33fF 
C361 tspc_1/Z2 VDD 0.91fF 
C362 tspc_1/Z1 VDD 0.41fF 
C363 tspc_0/Q VDD 1.95fF 
C364 nor_0/B VDD 4.86fF 
C365 tspc_0/a_630_n680# VDD 0.52fF 
C366 tspc_0/Z4 VDD 0.41fF 
C367 tspc_0/Z3 VDD 1.33fF 
C368 tspc_0/Z2 VDD 0.91fF 
C369 tspc_0/Z1 VDD 0.41fF 
C370 nor_0/A VDD 4.47fF 
C371 clk VDD 5.27fF 
C372 prescaler_0/nand_1/z1 VDD 0.20fF 
C373 prescaler_0/tspc_2/D VDD 1.94fF 
C374 and_0/OUT VDD 3.37fF 
C375 prescaler_0/nand_0/z1 VDD 0.20fF 
C376 vdd VDD 23.48fF 
C377 prescaler_0/tspc_1/Q VDD 1.91fF 
C378 prescaler_0/tspc_2/Q VDD 2.54fF 
C379 prescaler_0/tspc_2/a_630_n680# VDD 0.52fF 
C380 prescaler_0/tspc_2/Z4 VDD 0.41fF 
C381 prescaler_0/tspc_2/Z3 VDD 1.33fF 
C382 prescaler_0/tspc_2/Z2 VDD 0.91fF 
C383 prescaler_0/tspc_2/Z1 VDD 0.41fF 
C384 prescaler_0/tspc_2/a_740_n680# VDD 1.37fF 
C385 prescaler_0/tspc_1/a_630_n680# VDD 0.52fF 
C386 prescaler_0/tspc_1/Z4 VDD 0.41fF 
C387 prescaler_0/tspc_1/Z3 VDD 1.33fF 
C388 prescaler_0/tspc_1/Z2 VDD 0.91fF 
C389 prescaler_0/tspc_1/Z1 VDD 0.41fF 
C390 prescaler_0/m1_2700_2190# VDD 3.36fF 
C391 prescaler_0/tspc_0/a_630_n680# VDD 0.52fF 
C392 gnd VDD 21.02fF 
C393 prescaler_0/tspc_0/Z4 VDD 0.41fF 
C394 prescaler_0/Out VDD 3.22fF 
C395 prescaler_0/tspc_0/Z3 VDD 1.33fF 
C396 prescaler_0/tspc_0/Z2 VDD 0.91fF 
C397 prescaler_0/tspc_0/Z1 VDD 0.41fF 
C398 prescaler_0/tspc_0/D VDD 1.69fF 
C399 prescaler_0/tspc_0/a_740_n680# VDD 1.37fF 
C400 nor_1/Z1 VDD 0.58fF 
C401 mc2 VDD 3.39fF 
C402 nor_0/Z1 VDD 0.58fF 


.tran 0.1n 100n

.control
set hcopypscolor = 1
set color0 = white
set color1 = black

run

plot out+2 clk

.endc
.end