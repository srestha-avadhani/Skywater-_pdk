magic
tech sky130A
timestamp 1640700690
<< nwell >>
rect -55 -15 245 610
<< nmos >>
rect 20 -210 35 -110
rect 145 -210 160 -110
<< pmos >>
rect 20 10 35 460
rect 145 10 160 460
<< ndiff >>
rect -20 -130 20 -110
rect -20 -155 -15 -130
rect 10 -155 20 -130
rect -20 -175 20 -155
rect -20 -200 -15 -175
rect 10 -200 20 -175
rect -20 -210 20 -200
rect 35 -130 75 -110
rect 35 -155 45 -130
rect 70 -155 75 -130
rect 35 -175 75 -155
rect 35 -200 45 -175
rect 70 -200 75 -175
rect 35 -210 75 -200
rect 105 -130 145 -110
rect 105 -155 110 -130
rect 135 -155 145 -130
rect 105 -175 145 -155
rect 105 -200 110 -175
rect 135 -200 145 -175
rect 105 -210 145 -200
rect 160 -130 200 -110
rect 160 -155 170 -130
rect 195 -155 200 -130
rect 160 -175 200 -155
rect 160 -200 170 -175
rect 195 -200 200 -175
rect 160 -210 200 -200
<< pdiff >>
rect -20 450 20 460
rect -20 425 -15 450
rect 10 425 20 450
rect -20 405 20 425
rect -20 380 -15 405
rect 10 380 20 405
rect -20 360 20 380
rect -20 335 -15 360
rect 10 335 20 360
rect -20 315 20 335
rect -20 290 -15 315
rect 10 290 20 315
rect -20 270 20 290
rect -20 245 -15 270
rect 10 245 20 270
rect -20 225 20 245
rect -20 200 -15 225
rect 10 200 20 225
rect -20 180 20 200
rect -20 155 -15 180
rect 10 155 20 180
rect -20 135 20 155
rect -20 110 -15 135
rect 10 110 20 135
rect -20 90 20 110
rect -20 65 -15 90
rect 10 65 20 90
rect -20 45 20 65
rect -20 20 -15 45
rect 10 20 20 45
rect -20 10 20 20
rect 35 450 75 460
rect 35 425 45 450
rect 70 425 75 450
rect 35 405 75 425
rect 35 380 45 405
rect 70 380 75 405
rect 35 360 75 380
rect 35 335 45 360
rect 70 335 75 360
rect 35 315 75 335
rect 35 290 45 315
rect 70 290 75 315
rect 35 270 75 290
rect 35 245 45 270
rect 70 245 75 270
rect 35 225 75 245
rect 35 200 45 225
rect 70 200 75 225
rect 35 180 75 200
rect 35 155 45 180
rect 70 155 75 180
rect 35 135 75 155
rect 35 110 45 135
rect 70 110 75 135
rect 35 90 75 110
rect 35 65 45 90
rect 70 65 75 90
rect 35 45 75 65
rect 35 20 45 45
rect 70 20 75 45
rect 35 10 75 20
rect 105 450 145 460
rect 105 425 110 450
rect 135 425 145 450
rect 105 405 145 425
rect 105 380 110 405
rect 135 380 145 405
rect 105 360 145 380
rect 105 335 110 360
rect 135 335 145 360
rect 105 315 145 335
rect 105 290 110 315
rect 135 290 145 315
rect 105 270 145 290
rect 105 245 110 270
rect 135 245 145 270
rect 105 225 145 245
rect 105 200 110 225
rect 135 200 145 225
rect 105 180 145 200
rect 105 155 110 180
rect 135 155 145 180
rect 105 135 145 155
rect 105 110 110 135
rect 135 110 145 135
rect 105 90 145 110
rect 105 65 110 90
rect 135 65 145 90
rect 105 45 145 65
rect 105 20 110 45
rect 135 20 145 45
rect 105 10 145 20
rect 160 450 200 460
rect 160 425 170 450
rect 195 425 200 450
rect 160 405 200 425
rect 160 380 170 405
rect 195 380 200 405
rect 160 360 200 380
rect 160 335 170 360
rect 195 335 200 360
rect 160 315 200 335
rect 160 290 170 315
rect 195 290 200 315
rect 160 270 200 290
rect 160 245 170 270
rect 195 245 200 270
rect 160 225 200 245
rect 160 200 170 225
rect 195 200 200 225
rect 160 180 200 200
rect 160 155 170 180
rect 195 155 200 180
rect 160 135 200 155
rect 160 110 170 135
rect 195 110 200 135
rect 160 90 200 110
rect 160 65 170 90
rect 195 65 200 90
rect 160 45 200 65
rect 160 20 170 45
rect 195 20 200 45
rect 160 10 200 20
<< ndiffc >>
rect -15 -155 10 -130
rect -15 -200 10 -175
rect 45 -155 70 -130
rect 45 -200 70 -175
rect 110 -155 135 -130
rect 110 -200 135 -175
rect 170 -155 195 -130
rect 170 -200 195 -175
<< pdiffc >>
rect -15 425 10 450
rect -15 380 10 405
rect -15 335 10 360
rect -15 290 10 315
rect -15 245 10 270
rect -15 200 10 225
rect -15 155 10 180
rect -15 110 10 135
rect -15 65 10 90
rect -15 20 10 45
rect 45 425 70 450
rect 45 380 70 405
rect 45 335 70 360
rect 45 290 70 315
rect 45 245 70 270
rect 45 200 70 225
rect 45 155 70 180
rect 45 110 70 135
rect 45 65 70 90
rect 45 20 70 45
rect 110 425 135 450
rect 110 380 135 405
rect 110 335 135 360
rect 110 290 135 315
rect 110 245 135 270
rect 110 200 135 225
rect 110 155 135 180
rect 110 110 135 135
rect 110 65 135 90
rect 110 20 135 45
rect 170 425 195 450
rect 170 380 195 405
rect 170 335 195 360
rect 170 290 195 315
rect 170 245 195 270
rect 170 200 195 225
rect 170 155 195 180
rect 170 110 195 135
rect 170 65 195 90
rect 170 20 195 45
<< psubdiff >>
rect 230 -215 290 -155
<< nsubdiff >>
rect 95 540 145 590
<< poly >>
rect 20 460 35 480
rect 145 460 160 480
rect 20 -10 35 10
rect 145 -10 160 10
rect -20 -20 35 -10
rect -20 -40 -10 -20
rect 10 -40 35 -20
rect -20 -50 35 -40
rect 105 -20 160 -10
rect 105 -40 115 -20
rect 135 -40 160 -20
rect 105 -50 160 -40
rect 20 -110 35 -50
rect 145 -110 160 -50
rect 20 -225 35 -210
rect 145 -225 160 -210
<< polycont >>
rect -10 -40 10 -20
rect 115 -40 135 -20
<< locali >>
rect 90 535 150 595
rect 5 495 10 515
rect -15 460 10 495
rect -20 450 15 460
rect -20 425 -15 450
rect 10 425 15 450
rect -20 405 15 425
rect -20 380 -15 405
rect 10 380 15 405
rect -20 360 15 380
rect -20 335 -15 360
rect 10 335 15 360
rect -20 315 15 335
rect -20 290 -15 315
rect 10 290 15 315
rect -20 270 15 290
rect -20 245 -15 270
rect 10 245 15 270
rect -20 225 15 245
rect -20 200 -15 225
rect 10 200 15 225
rect -20 180 15 200
rect -20 155 -15 180
rect 10 155 15 180
rect -20 135 15 155
rect -20 110 -15 135
rect 10 110 15 135
rect -20 90 15 110
rect -20 65 -15 90
rect 10 65 15 90
rect -20 45 15 65
rect -20 20 -15 45
rect 10 20 15 45
rect -20 10 15 20
rect 40 450 75 460
rect 40 425 45 450
rect 70 425 75 450
rect 40 405 75 425
rect 40 380 45 405
rect 70 380 75 405
rect 40 360 75 380
rect 40 335 45 360
rect 70 335 75 360
rect 40 315 75 335
rect 40 290 45 315
rect 70 290 75 315
rect 40 270 75 290
rect 40 245 45 270
rect 70 245 75 270
rect 40 225 75 245
rect 105 450 140 460
rect 105 425 110 450
rect 135 425 140 450
rect 105 405 140 425
rect 105 380 110 405
rect 135 380 140 405
rect 105 360 140 380
rect 105 335 110 360
rect 135 335 140 360
rect 105 315 140 335
rect 105 290 110 315
rect 135 290 140 315
rect 105 270 140 290
rect 105 245 110 270
rect 135 245 140 270
rect 105 225 140 245
rect 40 200 45 225
rect 70 200 110 225
rect 135 200 140 225
rect 40 180 75 200
rect 40 155 45 180
rect 70 155 75 180
rect 40 135 75 155
rect 40 110 45 135
rect 70 110 75 135
rect 40 90 75 110
rect 40 65 45 90
rect 70 65 75 90
rect 40 45 75 65
rect 40 20 45 45
rect 70 20 75 45
rect 40 10 75 20
rect 105 180 140 200
rect 105 155 110 180
rect 135 155 140 180
rect 105 135 140 155
rect 105 110 110 135
rect 135 110 140 135
rect 105 90 140 110
rect 105 65 110 90
rect 135 65 140 90
rect 105 45 140 65
rect 105 20 110 45
rect 135 20 140 45
rect 105 10 140 20
rect 165 450 200 460
rect 165 425 170 450
rect 195 425 200 450
rect 165 405 200 425
rect 165 380 170 405
rect 195 380 200 405
rect 165 360 200 380
rect 165 335 170 360
rect 195 335 200 360
rect 165 315 200 335
rect 165 290 170 315
rect 195 290 200 315
rect 165 270 200 290
rect 165 245 170 270
rect 195 245 200 270
rect 165 225 200 245
rect 165 200 170 225
rect 195 200 200 225
rect 165 180 200 200
rect 165 155 170 180
rect 195 155 200 180
rect 165 135 200 155
rect 165 110 170 135
rect 195 110 200 135
rect 165 90 200 110
rect 165 65 170 90
rect 195 65 200 90
rect 165 45 200 65
rect 165 20 170 45
rect 195 20 200 45
rect 165 10 200 20
rect -20 -20 20 -10
rect -55 -40 -10 -20
rect 10 -40 20 -20
rect -20 -50 20 -40
rect 105 -20 145 -10
rect 105 -40 115 -20
rect 135 -40 145 -20
rect 105 -50 145 -40
rect 170 -70 195 10
rect 45 -90 245 -70
rect 45 -110 70 -90
rect 170 -110 195 -90
rect -20 -130 15 -110
rect -20 -155 -15 -130
rect 10 -155 15 -130
rect -20 -175 15 -155
rect -20 -200 -15 -175
rect 10 -200 15 -175
rect -20 -210 15 -200
rect 40 -130 75 -110
rect 40 -155 45 -130
rect 70 -155 75 -130
rect 40 -175 75 -155
rect 40 -200 45 -175
rect 70 -200 75 -175
rect 40 -210 75 -200
rect 105 -130 140 -110
rect 105 -155 110 -130
rect 135 -155 140 -130
rect 105 -175 140 -155
rect 105 -200 110 -175
rect 135 -200 140 -175
rect 105 -210 140 -200
rect 165 -130 200 -110
rect 165 -155 170 -130
rect 195 -155 200 -130
rect 165 -175 200 -155
rect 165 -200 170 -175
rect 195 -200 200 -175
rect 165 -210 200 -200
rect -15 -265 10 -210
rect 5 -285 10 -265
rect 110 -265 135 -210
rect 230 -215 290 -155
rect 130 -285 135 -265
<< viali >>
rect -15 495 5 515
rect 115 -40 135 -20
rect -15 -285 5 -265
rect 110 -285 130 -265
<< metal1 >>
rect -25 520 15 525
rect -25 490 -20 520
rect 10 490 15 520
rect -25 485 15 490
rect 105 -20 145 -10
rect 105 -40 115 -20
rect 135 -40 145 -20
rect 105 -50 145 -40
rect 115 -75 135 -50
rect -55 -90 135 -75
rect -25 -260 15 -255
rect -25 -290 -20 -260
rect 10 -290 15 -260
rect -25 -295 15 -290
rect 100 -260 140 -255
rect 100 -290 105 -260
rect 135 -290 140 -260
rect 100 -295 140 -290
<< via1 >>
rect -20 515 10 520
rect -20 495 -15 515
rect -15 495 5 515
rect 5 495 10 515
rect -20 490 10 495
rect -20 -265 10 -260
rect -20 -285 -15 -265
rect -15 -285 5 -265
rect 5 -285 10 -265
rect -20 -290 10 -285
rect 105 -265 135 -260
rect 105 -285 110 -265
rect 110 -285 130 -265
rect 130 -285 135 -265
rect 105 -290 135 -285
<< metal2 >>
rect -30 520 20 530
rect -30 490 -20 520
rect 10 490 20 520
rect -30 480 20 490
rect -30 -260 20 -250
rect -30 -290 -20 -260
rect 10 -290 20 -260
rect -30 -300 20 -290
rect 95 -260 145 -250
rect 95 -290 105 -260
rect 135 -290 145 -260
rect 95 -300 145 -290
<< via2 >>
rect -20 490 10 520
rect -20 -290 10 -260
rect 105 -290 135 -260
<< metal3 >>
rect -30 525 20 530
rect -30 485 -25 525
rect 15 485 20 525
rect -30 480 20 485
rect -30 -255 20 -250
rect -30 -295 -25 -255
rect 15 -295 20 -255
rect -30 -300 20 -295
rect 95 -255 145 -250
rect 95 -295 100 -255
rect 140 -295 145 -255
rect 95 -300 145 -295
<< via3 >>
rect -25 520 15 525
rect -25 490 -20 520
rect -20 490 10 520
rect 10 490 15 520
rect -25 485 15 490
rect -25 -260 15 -255
rect -25 -290 -20 -260
rect -20 -290 10 -260
rect 10 -290 15 -260
rect -25 -295 15 -290
rect 100 -260 140 -255
rect 100 -290 105 -260
rect 105 -290 135 -260
rect 135 -290 140 -260
rect 100 -295 140 -290
<< metal4 >>
rect -30 525 20 530
rect -55 495 -25 525
rect -30 485 -25 495
rect 15 495 245 525
rect 15 485 20 495
rect -30 480 20 485
rect -30 -255 20 -250
rect -30 -260 -25 -255
rect -55 -290 -25 -260
rect -30 -295 -25 -290
rect 15 -260 20 -255
rect 95 -255 145 -250
rect 95 -260 100 -255
rect 15 -290 100 -260
rect 15 -295 20 -290
rect -30 -300 20 -295
rect 95 -295 100 -290
rect 140 -260 145 -255
rect 140 -290 245 -260
rect 140 -295 145 -290
rect 95 -300 145 -295
<< labels >>
rlabel locali 110 565 110 565 1 vdd!
rlabel locali 265 -185 265 -185 1 gnd!
rlabel metal4 -55 -290 245 -260 1 GND
rlabel nwell -55 495 245 525 1 VDD
rlabel locali 75 200 105 225 1 Z1
rlabel locali 170 -90 245 -70 1 Out
rlabel locali -55 -40 10 -20 1 A
rlabel metal1 -55 -90 10 -75 1 B
<< end >>
