magic
tech sky130A
timestamp 1640777101
<< nwell >>
rect 0 580 1435 690
<< viali >>
rect 30 320 50 340
rect 1080 280 1100 300
rect 1435 280 1455 300
rect 30 -385 50 -365
<< metal1 >>
rect 20 345 60 350
rect 20 315 25 345
rect 55 315 60 345
rect 20 310 60 315
rect 1005 335 1050 350
rect 1200 335 1470 350
rect 1005 300 1020 335
rect 1070 300 1110 310
rect 1070 285 1080 300
rect 1020 280 1080 285
rect 1100 280 1110 300
rect 1020 270 1110 280
rect 1425 305 1465 310
rect 1425 275 1430 305
rect 1460 275 1465 305
rect 1425 270 1465 275
rect 1020 215 1035 270
rect 1020 200 1470 215
rect 20 -360 60 -355
rect 1020 -360 1035 200
rect 20 -390 25 -360
rect 55 -390 60 -360
rect 20 -395 60 -390
<< via1 >>
rect 25 340 55 345
rect 25 320 30 340
rect 30 320 50 340
rect 50 320 55 340
rect 25 315 55 320
rect 1430 300 1460 305
rect 1430 280 1435 300
rect 1435 280 1455 300
rect 1455 280 1460 300
rect 1430 275 1460 280
rect 25 -365 55 -360
rect 25 -385 30 -365
rect 30 -385 50 -365
rect 50 -385 55 -365
rect 25 -390 55 -385
<< metal2 >>
rect -115 395 0 410
rect 20 345 60 350
rect 20 315 25 345
rect 55 315 60 345
rect 20 310 60 315
rect 1420 305 1470 315
rect 1420 295 1430 305
rect 415 280 1430 295
rect 420 265 505 280
rect 1420 275 1430 280
rect 1460 275 1470 305
rect 1420 265 1470 275
rect 490 -310 505 265
rect 425 -325 505 -310
rect 15 -360 65 -350
rect 15 -390 25 -360
rect 55 -390 65 -360
rect 15 -400 65 -390
rect -115 -455 0 -440
<< via2 >>
rect 25 315 55 345
rect 25 -390 55 -360
<< metal3 >>
rect 15 350 65 355
rect 15 310 20 350
rect 60 310 65 350
rect 15 305 65 310
rect 15 -355 65 -350
rect 15 -395 20 -355
rect 60 -395 65 -355
rect 15 -400 65 -395
<< via3 >>
rect 20 345 60 350
rect 20 315 25 345
rect 25 315 55 345
rect 55 315 60 345
rect 20 310 60 315
rect 20 -360 60 -355
rect 20 -390 25 -360
rect 25 -390 55 -360
rect 55 -390 60 -360
rect 20 -395 60 -390
<< metal4 >>
rect -70 640 20 670
rect -70 350 -40 640
rect 15 350 65 355
rect -70 320 20 350
rect -70 -360 -40 320
rect 15 310 20 320
rect 60 310 65 350
rect 15 305 65 310
rect 10 -65 1020 20
rect 15 -355 65 -350
rect 15 -360 20 -355
rect -70 -390 20 -360
rect -70 -685 -40 -390
rect 15 -395 20 -390
rect 60 -395 65 -355
rect 15 -400 65 -395
rect -70 -715 20 -685
use and_pd  and_pd_0
timestamp 1640776259
transform 1 0 1100 0 1 395
box -120 -375 335 275
use tspc_r  tspc_r_1
timestamp 1640770827
transform 1 0 145 0 -1 -425
box -145 -380 875 305
use tspc_r  tspc_r_0
timestamp 1640770827
transform 1 0 145 0 1 380
box -145 -380 875 305
<< labels >>
rlabel nwell 980 600 1050 630 1 VDD
rlabel nwell 980 630 1020 640 1 VDD
rlabel space 985 50 1020 120 1 GND
rlabel space 985 85 1050 120 1 GND
rlabel metal4 10 -65 1020 20 1 GND
rlabel metal4 -70 -715 -40 670 1 VDD
rlabel metal2 -115 395 -70 410 1 REF
rlabel metal2 -115 -455 -70 -440 1 DIV
rlabel metal1 1415 335 1470 350 1 UP
rlabel metal1 1415 200 1470 215 1 DOWN
rlabel metal2 1435 280 1460 305 1 R
rlabel metal2 1140 280 1185 295 1 R
<< end >>
