magic
tech sky130A
timestamp 1640608660
<< nwell >>
rect -40 -10 300 290
<< nmos >>
rect 30 -225 45 -125
rect 155 -225 170 -125
<< pmos >>
rect 30 10 45 210
rect 155 10 170 210
<< ndiff >>
rect -10 -145 30 -125
rect -10 -170 -5 -145
rect 20 -170 30 -145
rect -10 -190 30 -170
rect -10 -215 -5 -190
rect 20 -215 30 -190
rect -10 -225 30 -215
rect 45 -145 85 -125
rect 45 -170 55 -145
rect 80 -170 85 -145
rect 45 -190 85 -170
rect 45 -215 55 -190
rect 80 -215 85 -190
rect 45 -225 85 -215
rect 115 -145 155 -125
rect 115 -170 120 -145
rect 145 -170 155 -145
rect 115 -190 155 -170
rect 115 -215 120 -190
rect 145 -215 155 -190
rect 115 -225 155 -215
rect 170 -145 210 -125
rect 170 -170 180 -145
rect 205 -170 210 -145
rect 170 -190 210 -170
rect 170 -215 180 -190
rect 205 -215 210 -190
rect 170 -225 210 -215
<< pdiff >>
rect -10 180 30 210
rect -10 155 -5 180
rect 20 155 30 180
rect -10 135 30 155
rect -10 110 -5 135
rect 20 110 30 135
rect -10 90 30 110
rect -10 65 -5 90
rect 20 65 30 90
rect -10 45 30 65
rect -10 20 -5 45
rect 20 20 30 45
rect -10 10 30 20
rect 45 180 85 210
rect 45 155 55 180
rect 80 155 85 180
rect 45 135 85 155
rect 45 110 55 135
rect 80 110 85 135
rect 45 90 85 110
rect 45 65 55 90
rect 80 65 85 90
rect 45 45 85 65
rect 45 20 55 45
rect 80 20 85 45
rect 45 10 85 20
rect 115 180 155 210
rect 115 155 120 180
rect 145 155 155 180
rect 115 135 155 155
rect 115 110 120 135
rect 145 110 155 135
rect 115 90 155 110
rect 115 65 120 90
rect 145 65 155 90
rect 115 45 155 65
rect 115 20 120 45
rect 145 20 155 45
rect 115 10 155 20
rect 170 180 210 210
rect 170 155 180 180
rect 205 155 210 180
rect 170 135 210 155
rect 170 110 180 135
rect 205 110 210 135
rect 170 90 210 110
rect 170 65 180 90
rect 205 65 210 90
rect 170 45 210 65
rect 170 20 180 45
rect 205 20 210 45
rect 170 10 210 20
<< ndiffc >>
rect -5 -170 20 -145
rect -5 -215 20 -190
rect 55 -170 80 -145
rect 55 -215 80 -190
rect 120 -170 145 -145
rect 120 -215 145 -190
rect 180 -170 205 -145
rect 180 -215 205 -190
<< pdiffc >>
rect -5 155 20 180
rect -5 110 20 135
rect -5 65 20 90
rect -5 20 20 45
rect 55 155 80 180
rect 55 110 80 135
rect 55 65 80 90
rect 55 20 80 45
rect 120 155 145 180
rect 120 110 145 135
rect 120 65 145 90
rect 120 20 145 45
rect 180 155 205 180
rect 180 110 205 135
rect 180 65 205 90
rect 180 20 205 45
<< psubdiff >>
rect 245 -265 290 -220
<< nsubdiff >>
rect 250 90 280 120
<< poly >>
rect 30 210 45 230
rect 155 210 170 230
rect 30 -75 45 10
rect 155 -75 170 10
rect 15 -85 55 -75
rect 15 -105 25 -85
rect 45 -105 55 -85
rect 15 -115 55 -105
rect 140 -85 180 -75
rect 140 -105 150 -85
rect 170 -105 180 -85
rect 140 -115 180 -105
rect 30 -125 45 -115
rect 155 -125 170 -115
rect 30 -245 45 -225
rect 155 -245 170 -225
<< polycont >>
rect 25 -105 45 -85
rect 150 -105 170 -85
<< locali >>
rect -5 210 15 250
rect 120 210 140 250
rect -10 180 25 210
rect -10 155 -5 180
rect 20 155 25 180
rect -10 135 25 155
rect -10 110 -5 135
rect 20 110 25 135
rect -10 90 25 110
rect -10 65 -5 90
rect 20 65 25 90
rect -10 45 25 65
rect -10 20 -5 45
rect 20 20 25 45
rect -10 10 25 20
rect 50 180 85 210
rect 50 155 55 180
rect 80 155 85 180
rect 50 135 85 155
rect 50 110 55 135
rect 80 110 85 135
rect 50 90 85 110
rect 50 65 55 90
rect 80 65 85 90
rect 50 45 85 65
rect 50 20 55 45
rect 80 20 85 45
rect 50 10 85 20
rect 115 180 150 210
rect 115 155 120 180
rect 145 155 150 180
rect 115 135 150 155
rect 115 110 120 135
rect 145 110 150 135
rect 115 90 150 110
rect 115 65 120 90
rect 145 65 150 90
rect 115 45 150 65
rect 115 20 120 45
rect 145 20 150 45
rect 115 10 150 20
rect 175 180 210 210
rect 175 155 180 180
rect 205 155 210 180
rect 175 135 210 155
rect 175 110 180 135
rect 205 110 210 135
rect 175 90 210 110
rect 175 65 180 90
rect 205 65 210 90
rect 245 85 285 125
rect 175 45 210 65
rect 175 20 180 45
rect 205 20 210 45
rect 175 10 210 20
rect 60 -15 80 10
rect 185 -15 205 10
rect 60 -40 300 -15
rect 15 -85 55 -65
rect 140 -85 180 -65
rect -25 -105 25 -85
rect 45 -105 55 -85
rect 100 -105 150 -85
rect 170 -105 180 -85
rect -10 -145 25 -125
rect -10 -170 -5 -145
rect 20 -170 25 -145
rect -10 -190 25 -170
rect -10 -215 -5 -190
rect 20 -215 25 -190
rect -10 -225 25 -215
rect 50 -145 85 -125
rect 115 -145 150 -125
rect 50 -170 55 -145
rect 80 -170 120 -145
rect 145 -170 150 -145
rect 50 -190 85 -170
rect 50 -215 55 -190
rect 80 -215 85 -190
rect 50 -225 85 -215
rect 115 -190 150 -170
rect 115 -215 120 -190
rect 145 -215 150 -190
rect 115 -225 150 -215
rect 175 -145 210 -125
rect 175 -170 180 -145
rect 205 -150 210 -145
rect 230 -150 250 -40
rect 205 -170 250 -150
rect 175 -190 210 -170
rect 175 -215 180 -190
rect 205 -215 210 -190
rect 175 -225 210 -215
rect -5 -275 20 -225
rect 240 -270 295 -215
rect 15 -295 20 -275
<< viali >>
rect -5 250 15 270
rect 120 250 140 270
rect 150 -105 170 -85
rect -5 -295 15 -275
<< metal1 >>
rect -15 275 25 280
rect -15 245 -10 275
rect 20 245 25 275
rect 110 275 150 280
rect 110 245 115 275
rect 145 245 150 275
rect -25 -60 170 -45
rect 155 -75 170 -60
rect 140 -85 180 -75
rect 140 -105 150 -85
rect 170 -105 180 -85
rect 140 -115 180 -105
rect -15 -270 25 -265
rect -15 -300 -10 -270
rect 20 -300 25 -270
<< via1 >>
rect -10 270 20 275
rect -10 250 -5 270
rect -5 250 15 270
rect 15 250 20 270
rect -10 245 20 250
rect 115 270 145 275
rect 115 250 120 270
rect 120 250 140 270
rect 140 250 145 270
rect 115 245 145 250
rect -10 -275 20 -270
rect -10 -295 -5 -275
rect -5 -295 15 -275
rect 15 -295 20 -275
rect -10 -300 20 -295
<< metal2 >>
rect -15 275 25 280
rect -15 245 -10 275
rect 20 245 25 275
rect -15 240 25 245
rect 110 275 150 280
rect 110 245 115 275
rect 145 245 150 275
rect 110 240 150 245
rect -15 -270 25 -265
rect -15 -300 -10 -270
rect 20 -300 25 -270
rect -15 -305 25 -300
<< via2 >>
rect -10 245 20 275
rect 115 245 145 275
rect -10 -300 20 -270
<< metal3 >>
rect -20 280 30 285
rect -20 245 -10 280
rect 25 245 30 280
rect -20 235 30 245
rect 105 280 155 285
rect 105 245 115 280
rect 150 245 155 280
rect 105 235 155 245
rect -20 -265 30 -260
rect -20 -305 -15 -265
rect 25 -305 30 -265
rect -20 -310 30 -305
<< via3 >>
rect -10 275 25 280
rect -10 245 20 275
rect 20 245 25 275
rect 115 275 150 280
rect 115 245 145 275
rect 145 245 150 275
rect -15 -270 25 -265
rect -15 -300 -10 -270
rect -10 -300 20 -270
rect 20 -300 25 -270
rect -15 -305 25 -300
<< metal4 >>
rect -40 280 275 290
rect -40 260 -10 280
rect -20 245 -10 260
rect 25 260 115 280
rect 25 245 30 260
rect -20 235 30 245
rect 105 245 115 260
rect 150 260 275 280
rect 150 245 155 260
rect 105 235 155 245
rect -20 -265 30 -260
rect -20 -305 -15 -265
rect 25 -280 30 -265
rect 25 -305 275 -280
rect -20 -310 275 -305
<< labels >>
rlabel locali 60 -40 250 -15 1 OUT
rlabel space 100 -105 170 -85 1 B
rlabel locali -25 -105 45 -85 1 A
rlabel locali 265 100 265 100 1 vdd!
rlabel locali 265 -245 265 -245 1 gnd!
rlabel nwell -40 260 275 290 1 VDD
rlabel metal4 -20 -310 275 -280 1 GND
rlabel locali 55 -170 145 -145 1 z1
<< end >>
